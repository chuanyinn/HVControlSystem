* AD5686R SPICE Macro-model
* Description: Digital to Analog Converter
* Revision History:
*   Rev.1.0 Nov 2016
* Copyright 2016 by Analog Devices, Inc.
*
* Refer to http://www.analog.com/Analog_Root/static/techSupport/designTools/spiceModels/license/spice_general.html
* for License Statement. Use of this model indicates your acceptance
* of the terms and provisions in the License Staement.
*
* BEGIN Notes:
*
* The serial interface (SYNC, SCLK, SDIN, SDO) and the LDAC pin have been replaced with a simple parallel interface in this model.
* This makes it easier to load input data during simulation.
* Parallel interface description:
*   IN[0:15]   16 bit parallel input data
*   STROBE     Data on IN[0:16] is loaded into the input register on the rising edge of STROBE
*   DACLoad    The DAC Output is updated on the rising  edge of DAC_LOAD
*   CH_*       When high the corresponding channel will be updated on the rising edge of DAC_LOAD

* Not modeled: Serial Interface functionality and timing, SCLK pin, SYNC pin, SDIN pin, SDO pin, LDAC pin, 
*              daisy chain and readback modes, Software functions, noise, Turn On/Turn Off time 
*
* Parameters modeled include:
*    Slew Rate, Settling time, Resolution, Zero Code Error, Offset Error, Gain Error
*    Crosstalk, Short Circuit current, Quiescent supply currents,
*    RESETB and RSTSEL pin functionality, GAIN pin functionality
* 
* This model will not run in Multisim.
*  
* END Notes
* 
.param vscale={1/10000}
.param cscale=1e-5
.param rscale={1/cscale}
.PARAM ref_val=2.5
+ PwrOn=0
+ Ref_Sel = 0
+ PSRR_EN = 1
+ gain_error = 0
+ zero_code_error = 0.4m
+ dnl_en = 1
+ offs_error = 0.1m
+ crosstalk_en = 1
+ Dc_gain = 899999999.77
+ Freq3dB = 0.1
+ slewrate = 0.8
+ Rout = 23.717
.SUBCKT AD5686R CH_A CH_B CH_C CH_D DACLoad
+  GAIN GND IN0 IN1 IN2 IN3 IN4 IN5 IN6 IN7 IN8 IN9 IN10 IN11 IN12 IN13 IN14 IN15
+  RESETB RSTSEL STROBE VDD VLOGIC VOUTA VOUTB VOUTC VOUTD VREF 
X_dr9 CH_C DACLOAD_EDGE_TRIGER_INT IN_REG_OUT DAC_C 
+  RST_MIDCODE_INT RST_ZERO_INT DAC_Reg  
R_R8         N1698899 OUTA_INT  1m   
X_c11 VOUTB_INT VOUTB Current_Limit_ckt  
C_C9         OUTD_INT 0  1n  IC=0  
C_C7         OUTB_INT 0  1n  IC=0  
X_dr8 CH_B DACLOAD_EDGE_TRIGER_INT IN_REG_OUT DAC_B 
+ RST_MIDCODE_INT RST_ZERO_INT DAC_Reg  
X_dr10 CH_D DACLOAD_EDGE_TRIGER_INT IN_REG_OUT DAC_D 
+ RST_MIDCODE_INT RST_ZERO_INT DAC_Reg  
C_C6         OUTA_INT 0  1n IC=0   
C_C8         OUTC_INT 0  1n IC=0
X_dac1 DAC_A N1698899 DAC_REF DAC  
R_R11         N1593807 OUTD_INT  1m   
X_c1 VOUTA_INT VOUTA Current_Limit_ckt  
R_R9         N1698994 OUTB_INT  1m   
X_c12 VOUTC_INT VOUTC Current_Limit_ckt  
X_dr1 CH_A DACLOAD_EDGE_TRIGER_INT  IN_REG_OUT DAC_A 
+ RST_MIDCODE_INT RST_ZERO_INT DAC_Reg  
X_c13 VOUTD_INT VOUTD Current_Limit_ckt PARAMS: ILIMITN=40m ILIMITP=40m
R_R10         N1593799 OUTC_INT  1m   
E_ABM7         INT_REF_SEL 0 VALUE { 1-V(REF_SEL)    }
*.IC         V(VREF )=2.5
X_dig1 DACLOAD DACLOAD_EDGE_TRIGER_INT GAIN GAIN_FACTOR_INT
+  RESETB RST_MIDCODE_INT RST_ZERO_INT RSTSEL STROBE STROBE_EDGE_TRIGER_INT
+  VLOGIC_INT Internal_Logic  
V_V75         VREF_INT 0 {ref_val}
E_ABM11         DAC_REF 0 VALUE { if(Ref_Sel>0.8,V(VREF),V(VREF_INT))    }
X_Ref1 INTERNAL_REF VREF_INT INTERNAL_REF VDD_INT Reference_Buffer   
X_power1 GND REF_SEL VDD VDD_INT VLOGIC VLOGIC_INT Current_Model  
V_V74         REF_SEL 0 {Ref_Sel}
X_In1 IN0 IN1 IN2 IN3 IN4 IN5 IN6 IN7 IN8 IN9 IN10 IN11 IN12 IN13 IN14 IN15
+  IN_REG_OUT RST_MIDCODE_INT RST_ZERO_INT STROBE_EDGE_TRIGER_INT
+  InputReg_Bin_Dec  
X_s2 INTERNAL_REF VREF INT_REF_SEL switch_ideal  
*.IC         V(INTERNAL_REF )=2.5
X_ps1 0 PSRR_ADD VDD_INT DC_PSRR 
X_limit1 VDD Voltage_CLamp PARAMS: HIGH=5.51 LOW=2.7
X_limit2 VLOGIC Voltage_CLamp PARAMS: HIGH=5.51 LOW=1.8
X_dac11 DAC_B N1698994 DAC_REF DAC  
X_dac12 DAC_C N1593799 DAC_REF DAC  
X_dac13 DAC_D N1593807 DAC_REF DAC  
X_op2 N1789987 VOUTA_CHNL VOUTA_INT VDD_INT 0 opamp_parameterised  
X_Top1_S3    GAIN_FACTOR_INT 0 N1789987 0 AD5560_Top_Top1_S3 
R_R12         N1789987 VOUTA_INT  10k   
X_ctalk1 N1790473 CH_B CH_C CH_D GAIN_FACTOR_INT
+  VOUTB_INT VOUTC_INT VOUTD_INT Crosstalk  
E_ABM1         VOUTA_CHNL 0 VALUE { ( V(N1790473)  
+ +V(OUTA_INT)  
+ +V(PSRR_ADD))  }
X_Top1_S4    GAIN_FACTOR_INT 0 N1791678 0 AD5560_Top_Top1_S4 
X_op8 N1791678 VOUTB_CHNL VOUTB_INT VDD_INT 0 opamp_parameterised  
R_R13         N1791678 VOUTB_INT  10k   
X_ctalk2 N1792173 CH_A CH_C CH_D GAIN_FACTOR_INT
+  VOUTA_INT VOUTC_INT VOUTD_INT Crosstalk  
E_ABM8         VOUTB_CHNL 0 VALUE { ( V(N1792173)  
+ +V(OUTB_INT)  
+ +V(PSRR_ADD))  }
X_Top1_S5    GAIN_FACTOR_INT 0 N1793310 0 AD5560_Top_Top1_S5 
X_op9 N1793310 VOUTC_CHNL VOUTC_INT VDD_INT 0 opamp_parameterised  
R_R14         N1793310 VOUTC_INT  10k   
E_ABM9         VOUTC_CHNL 0 VALUE { ( V(N1793792)  
+ +V(OUTC_INT)  
+ +V(PSRR_ADD))  }
X_ctalk3 N1793792 CH_B CH_A CH_D GAIN_FACTOR_INT
+  VOUTB_INT VOUTA_INT VOUTD_INT Crosstalk  
R_R15         N1794947 VOUTD_INT  10k   
X_Top1_S6    GAIN_FACTOR_INT 0 N1794947 0 AD5560_Top_Top1_S6 
X_op10 N1794947 VOUTD_CHNL VOUTD_INT VDD_INT 0 opamp_parameterised  
E_ABM10         VOUTD_CHNL 0 VALUE { ( V(N1795428)  
+ +V(OUTD_INT)  
+ +V(PSRR_ADD))  }
X_ctalk4 N1795428 CH_B CH_C CH_A GAIN_FACTOR_INT
+  VOUTB_INT VOUTC_INT VOUTA_INT Crosstalk 
X_limit3 VOUTA Voltage_CLamp PARAMS: HIGH=5.5001 LOW=0
X_limit4 VOUTB Voltage_CLamp PARAMS: HIGH=5.5001 LOW=0
X_limit5 VOUTC Voltage_CLamp PARAMS: HIGH=5.5001 LOW=0
X_limit6 VOUTD Voltage_CLamp PARAMS: HIGH=5.5001 LOW=0 
.ENDS AD5686R
*$ Top Level Main Ends Here *$
.SUBCKT Crosstalk crosstalk_out en1 en2 en3 gain_factor out1 out2 out3 
V_V1         CROSSTALK_EN 0 {crosstalk_en}
E_TABLE1         N887992 0 TABLE {V(OUTPUT_CHANGE)} 0V           0V  
+ 0.5V           4e-7V  
+ 1V           8e-7V  
+ 1.5V           1.2e-6V  
+ 2.5V           2e-6V
E_ABM2         CROSSTALK_OUT 0 VALUE { if(V(CROSSTALK_EN)>0.5,V(N887992),0)    
+  }
E_ABM1         OUTPUT_CHANGE 0 VALUE {
+  (V(OUT1)*V(EN1))+(V(OUT2)*V(EN2))+(V(OUT3)*V(EN3))    }
.ENDS Crosstalk 
*$ 
.subckt opamp_parameterised INM INP out VDD VSS
R1 R1_P N1796906 8k
R_R4 0 N1763459  { (1*slewrate*1e6) /(6.28*Freq3dB) }
R_R13 N1797044 0  1
R_R14 N1796906 0 {1meg-8000}
R_R9 OUT 0  {Rout}
V_V7 K 0  { (Dc_gain*Freq3dB*6.28) / (slewrate*1e6) }


C_C10 0 N1797044  61.826n ; IC 0  


C_C11 R1_P 0  20u ; IC 0  

G_ABM2I3 0 N1763459  VALUE { LIMIT((V(K)*V(inp,inm)),-125,125) }
G1 N1797044 0 N1796906 0 -1 
G2 N1796906 0 N1763459 0 {-1/(1meg-8000)} 
G3 OUT 0 N1797044 0 {-1/ROUT} 


C_C8 0 N1763459  {1/ (slewrate*1e6) } ; IC 0  

.ends opamp_parameterised

*$ 
.SUBCKT Voltage_CLamp limit_node PARAMS: HIGH=5.5 LOW=2.7
V_V187         N1409984 0 {high}
V_V188         N1409988 0 {low}
X_U98         LIMIT_NODE N1409984 DIODE
X_U99         N1409988 LIMIT_NODE DIODE
.ENDS Voltage_CLamp 
*$ 
.SUBCKT DC_PSRR GND PSRR_ADD VDD 
E_ABM3         PSRR_ADD 0 VALUE { if(V(PSRR_EN)>0.5,V(PSRR_INT),0)    }
V_V1         PSRR_EN 0 {PSRR_EN}
E_TABLE1         PSRR_INT 0 TABLE {V(VDD)} 0V        0mV  
+ 1.8V        0mV  
+ 2.7V       0mV  
+ 4.5V     -0.075mV  
+ 5.5V      0.075mV
.ENDS DC_PSRR 
*$ 
.SUBCKT switch_ideal in out Vth  
X_Top1_s2_S1    VTH 0 OUT IN switch_ideal_Top1_s2_S1 
.ENDS switch_ideal 
*$


.SUBCKT InputReg_Bin_Dec IN0 IN1 IN2 IN3 IN4 IN5 IN6 IN7 IN8 IN9 IN10 IN11 IN12
+  IN13 IN14 IN15 Input_Reg_out rst_midcode rst_zero strobe  
X_b1 DEC_OUT IN0_INT IN1_INT IN2_INT IN3_INT IN4_INT IN5_INT IN6_INT IN7_INT
+  IN8_INT IN9_INT IN10_INT IN11_INT IN12_INT IN13_INT IN14_INT IN15_INT BintoDec
+   
R_R16         N1713111 INT_OUT  {10m*rscale}   
E_ABM16         N1713111 0 VALUE { IF(V(STROBE)>.9,V(DEC_OUT)*vscale,V(INT_OUT))     }
E_E1         INPUT_REG_OUT 0 INT_OUT 0 {1/vscale}
C_C17         0 INT_OUT  {1n*cscale} IC=0   
E_ABM6         N1720992 0 VALUE { IF(V(RST_MIDCODE)>.9,32768*vscale,V(INT_OUT))     }
R_R2         INT_OUT N1721034  {1m*rscale}
E_ABM7         N1721034 0 VALUE { IF(V(RST_ZERO)>.9,0,V(INT_OUT))     }
R_R4         INT_OUT N1720992  {1m*rscale}
E_ABM64         IN0_INT 0 VALUE { if(V(IN0)>0.5,1,0)    }
E_ABM65         IN1_INT 0 VALUE { if(V(IN1)>0.5,1,0)    }
E_ABM66         IN2_INT 0 VALUE { if(V(IN2)>0.5,1,0)    }
E_ABM67         IN3_INT 0 VALUE { if(V(IN3)>0.5,1,0)    }
E_ABM68         IN4_INT 0 VALUE { if(V(IN4)>0.5,1,0)    }
E_ABM69         IN5_INT 0 VALUE { if(V(IN5)>0.5,1,0)    }
E_ABM70         IN6_INT 0 VALUE { if(V(IN6)>0.5,1,0)    }
E_ABM71         IN7_INT 0 VALUE { if(V(IN7)>0.5,1,0)    }
E_ABM72         IN8_INT 0 VALUE { if(V(IN8)>0.5,1,0)    }
E_ABM73         IN9_INT 0 VALUE { if(V(IN9)>0.5,1,0)    }
E_ABM74         IN10_INT 0 VALUE { if(V(IN10)>0.5,1,0)    }
E_ABM75         IN11_INT 0 VALUE { if(V(IN11)>0.5,1,0)    }
E_ABM76         IN12_INT 0 VALUE { if(V(IN12)>0.5,1,0)    }
E_ABM77         IN13_INT 0 VALUE { if(V(IN13)>0.5,1,0)    }
E_ABM78         IN14_INT 0 VALUE { if(V(IN14)>0.5,1,0)    }
E_ABM79         IN15_INT 0 VALUE { if(V(IN15)>0.5,1,0)    }
.ENDS InputReg_Bin_Dec 
*$ 
.SUBCKT BintoDec dec_out InReg_out0 InReg_out1 InReg_out2 InReg_out3 InReg_out4
+  InReg_out5 InReg_out6 InReg_out7 InReg_out8 InReg_out9 InReg_out10 InReg_out11
+  InReg_out12 InReg_out13 InReg_out14 InReg_out15  
E_ABM1         OUT_1 0 VALUE {
+  ((V(INREG_OUT0)*1)+(V(INREG_OUT1)*PWR(2,1))+(V(INREG_OUT2)*PWR(2,2))  
+ +(V(INREG_OUT3)*PWR(2,3))+(V(INREG_OUT4)*PWR(2,4))+(V(INREG_OUT5)*PWR(2,5)) 
+  
+ +(V(INREG_OUT6)*PWR(2,6))+(V(INREG_OUT7)*PWR(2,7))+(V(INREG_OUT8)*PWR(2,8)) 
+  
+
+  +(V(INREG_OUT9)*PWR(2,9))+(V(INREG_OUT10)*PWR(2,10))+(V(INREG_OUT11)*PWR(2,11)))
+  }
E_ABM6         OUT_2 0 VALUE {
+  ((V(INREG_OUT12)*PWR(2,12))+(V(INREG_OUT13)*PWR(2,13))+(V(INREG_OUT14)*PWR(2,14))
+   
+ +(V(INREG_OUT15)*PWR(2,15)))   }
E_ABM7         DEC_OUT 0 VALUE { V(OUT_1)+V(OUT_2)    }
.ENDS BintoDec 
*$ 
.SUBCKT Current_Model GND REF_SEL VDD VDD_INT VLOGIC VLOGIC_INT  
E_E2         VLOGIC_INT GND VLOGIC GND 1
G_ABMI5         VLOGIC GND VALUE { 3u    }
E_E1         VDD_INT GND VDD GND 1
G_ABMI4         VDD GND VALUE { if(V(REF_SEL)<0.2,1.1m,0.59m)    }
.ENDS Current_Model 
*$ 


.subckt Reference_Buffer inm inp OUT VDD
R_R1 N1807677 0 {1-14m}
R_R2 OUT 0  3900
R1 R1_P N1807577 8k
R_R3 N1808025 N1807813  1
R2 R2_P N1807677 14m


R3 N1808025 0 1meg

R_R5 N1807577 0 {1Meg-8000}
R_R6 0 N1807673  { (1*1e6) / (6.28*0.1) }
V_V1 K 0  { 899999999*0.1*6.28 / (1*1e6) }


L_L4 N1808025 0  28u ;IC 0  

C_C11 R1_P 0 20u  


C_C12 R2_P 0  0.002 ;IC 2.5  

G_ABM2I3 0 N1807673 VALUE = { LIMIT((V(K)*V(INP,INM)),-1000,1000) }
G_G4 N1807813 0 N1807673 0  -1
G1 N1807577 0 N1807813 0 {-1/(1meg-8000)} 
G2 N1807677 0 N1807577 0 {-1/(1-14m)} 
G3 OUT 0 N1807677 0 {-1/3900} 


C_C8 0 N1807673  {1/ (1*1e6) } ;IC 2.5  

.ends Reference_Buffer



*$ 
.SUBCKT Internal_Logic DACLoad DACLoad_edge_triger GAIN gain_factor
+ RESETb rst_midcode rst_zero RSTSEL strobe strobe_edge_triger
+  VLOGIC  
X_U32         STROBE N1581148 INV_DELAY_SAN PARAMS: VDD=1 VSS=0 VTH=0.5
+  DELAY=16n
E_ABM1         RST_ZERO_INT 0 VALUE { if(V(RESETB)<0.1 & V(RSTSEL)<0.9,1,0)   
+  }
E_ABM2         RST_MIDCODE_INT 0 VALUE { if(V(RESETB)<0.1 & V(RSTSEL)>0.9,1,0) 
+    }
X_U36         RST_MIDCODE_INT N1585905 RST_MIDCODE AND2_SAN PARAMS:  VDD=1
+  VSS=0 VTH=0.5 DELAY=1e-11 
X_U35         RST_MIDCODE_INT N1585905 INV_DELAY_SAN PARAMS: VDD=1 VSS=0
+  VTH=0.5 DELAY=20n
X_U33         DACLOAD N1581384 N1581388 AND2_SAN PARAMS:  VDD=1
+  VSS=0 VTH=0.5 DELAY=1e-12 
X_U34         DACLOAD N1581384 INV_DELAY_SAN PARAMS: VDD=1 VSS=0 VTH=0.5
+  DELAY=15n
E_ABM8         GAIN_FACTOR 0 VALUE { if(V(GAIN)>0.9,2,1)    }
X_U1         STROBE N1581148 STROBE_EDGE_TRIGER AND2_SAN PARAMS:  VDD=1 VSS=0
+  VTH=0.5 DELAY=1e-12 
X_U38         RST_ZERO_INT N1750861 RST_ZERO AND2_SAN PARAMS:  VDD=1 VSS=0
+  VTH=0.5 DELAY=1e-12 
X_U37         RST_ZERO_INT N1750861 INV_DELAY_SAN PARAMS: VDD=1 VSS=0 VTH=0.5
+  DELAY=20n
X_U39         N1581388 RESETB DACLOAD_EDGE_TRIGER AND2_SAN PARAMS:  VDD=1 VSS=0
+  VTH=0.5 DELAY=1e-11
.ENDS Internal_Logic 
*$ 
.SUBCKT DAC code dacout Vref  
V_V2         GAIN_ERROR_LSB 0 {gain_error/(2**16-1)}
E_ABM1         DACOUT_INT 0 VALUE { V(LSB)*V(CODE)    }
X_U1         DNL_ERR CODE N887486 INL_ADD
E_ABM2         DC_ERROR 0 VALUE { offs_error+zero_code_error    }
E_ABM5         LSB 0 VALUE { (V(VREF)/(2**16))+V(GAIN_ERROR_LSB)    }
E_ABM4         DACOUT_WD_ERR 0 VALUE { ( V(DNL_ERR)  
+ +V(DAC_WD_DC_ERR) )   }
V_V1         N887486 0 {dnl_en}
E_ABM3         DAC_WD_DC_ERR 0 VALUE { ( V(DC_ERROR)  
+ +V(DACOUT_INT) )   }
E_ABM6         DACOUT 0 VALUE { LIMIT(V(DACOUT_WD_ERR),0,2.5)    }
.ENDS DAC 
*$ 
.SUBCKT Current_Limit_ckt I_in I_out PARAMS: ILIMITN=40M ILIMITP=40M
X_U22         N1248164 I_IN DIODE
I_I6         I_IN N1248164 DC {ilimitp}  
I_I7         I_OUT N1248164 DC {ilimitn}  
X_U21         N1248164 I_OUT DIODE
.ENDS Current_Limit_ckt 
*$ 
.SUBCKT DAC_Reg DAC_en DAC_load DACReg_in DACReg_out 
+  rst_midcode rst_zero  
R_R1         N1546964 INT_OUT  {1m*rscale}
C_C1         INT_OUT 0 {1n*cscale} IC={0+(PwrOn*32768)}  
E_E16         DACREG_OUT 0 INT_OUT 0 {1/vscale}
E_ABM1         N1546964 0 VALUE { IF(V(DAC_LOAD)>.9 & V(DAC_EN)>.9,V(DACReg_in)*vscale,V(INT_OUT))     }
E_ABM6         N1680667 0 VALUE { IF(V(RST_MIDCODE)>.9,32768*vscale,V(INT_OUT))     }
R_R4         INT_OUT N1680667  {1m*rscale}   
R_R2         INT_OUT N1720858  {1m*rscale}   
E_ABM7         N1720858 0 VALUE { IF(V(RST_ZERO)>.9,0,V(INT_OUT))     }
.ENDS DAC_Reg 
*$
.subckt AD5560_Top_Top1_S3 1 2 3 4  
S_S3         3 4 1 2 _S3
RS_S3         1 2 1G
.MODEL         _S3 VSWITCH Roff=1e10 Ron=10k Voff=1.3 Von=1.5
.ends AD5560_Top_Top1_S3
*$
.subckt AD5560_Top_Top1_S4 1 2 3 4  
S_S4         3 4 1 2 _S4
RS_S4         1 2 1G
.MODEL         _S4 VSWITCH Roff=1e10 Ron=10k Voff=1.3 Von=1.5
.ends AD5560_Top_Top1_S4
*$
.subckt AD5560_Top_Top1_S5 1 2 3 4  
S_S5         3 4 1 2 _S5
RS_S5         1 2 1G
.MODEL         _S5 VSWITCH Roff=1e10 Ron=10k Voff=1.3 Von=1.5
.ends AD5560_Top_Top1_S5
*$
.subckt AD5560_Top_Top1_S6 1 2 3 4  
S_S6         3 4 1 2 _S6
RS_S6         1 2 1G
.MODEL         _S6 VSWITCH Roff=1e10 Ron=10k Voff=1.3 Von=1.5
.ends AD5560_Top_Top1_S6
*$
.subckt switch_ideal_Top1_s2_S1 1 2 3 4  
S_S1         3 4 1 2 _S1
RS_S1         1 2 1G
.MODEL         _S1 VSWITCH Roff=1e10 Ron=1m Voff=0.45V Von=0.55V
.ends switch_ideal_Top1_s2_S1
*$
******************************* Other Subckts Used In Design ************************************
*$
.SUBCKT AND2_SAN IN1 IN2 OUT PARAMS:VDD=5 VSS=0 VTH=2.5 DELAY = 1p 
E1 OUT1 0 VALUE={if(V(IN1)>{VTH}&V(IN2)>{VTH},{VDD},{VSS})}
R1 OUT1 OUT2 {{DELAY}*1E12}
C1 OUT2 0 1.443p
E2 OUT 0 VALUE={IF(V(OUT2)>{VTH},{VDD},{VSS})}
.ENDS AND2_SAN
*$
.SUBCKT AND3_SAN IN1 IN2 IN3 OUT PARAMS:VDD=5 VSS=0 VTH=2.5 DELAY = 1N
E3 OUT1 0 VALUE={if(V(IN1)>{VTH}&V(IN2)>{VTH}&V(IN3)>{VTH},{VDD},{VSS})}
R3 OUT1 OUT {{DELAY}*1E9}
C3 OUT 0 1.443n
.ENDS AND3_SAN
*$
.SUBCKT AND4_SAN IN1 IN2 IN3 IN4 OUT PARAMS:VDD=5 VSS=0 VTH=2.5 DELAY=1n
E4 OUT1 0 VALUE={if(V(IN1)>{VTH}&V(IN2)>{VTH}&V(IN3)>{VTH}&V(IN4)>{VTH},{VDD},0)}
R4 OUT1 OUT {{DELAY}*1E9}
C4 OUT 0 1.443n
.ENDS AND4_SAN 
*$
*WITH DELAY
.SUBCKT BUF_DELAY_SAN IN OUT PARAMS: VDD=5 VSS=0 DELAY=1p VTH = 2.5
E1 OUT1 0 VALUE = {IF(V(IN)>{VTH},{VDD},{VSS})}
R1 OUT1 OUT2 {{DELAY}*1E12}
C1 OUT2 0 1.443p
E2 OUT 0 VALUE={IF(V(OUT2)>{VTH},{VDD},{VSS})}
.ENDS BUF_DELAY_SAN 
*DIODE
*$
.SUBCKT DIODE 1 2 
D1 1 2 ideal
.model ideal D n=1m is=1e-15 tt=1f rs=1n
.ENDS DIODE
*$
*WITH DELAY
.SUBCKT INV_DELAY_SAN IN OUT PARAMS: VDD=5 VSS=0 VTH=2.5 DELAY=1p
E1 OUT1 0 VALUE={IF(V(IN)>{VTH},{VSS},{VDD})}
R1 OUT1 OUT2 {{DELAY}*1E12}
C1 OUT2 0 1.443p
E2 OUT 0 VALUE={IF(V(OUT2)>{VTH},{VDD},{VSS})}
.ENDS INV_DELAY_SAN
*$
.SUBCKT NAND2_SAN IN1 IN2 OUT PARAMS:VDD=5 VSS=0 VTH=2.5 DELAY=1n
E3 OUT1 0 VALUE={if(V(IN1)>{VTH}&V(IN2)>{VTH},0,{VDD})}
R3 OUT1 OUT {{DELAY}*1E9}
C3 OUT 0 1.443n
.ENDS NAND2_SAN
*$
.SUBCKT NAND3_SAN IN1 IN2 IN3 OUT PARAMS:VDD=5 VSS=0 VTH=2.5 DELAY=1n
E3 OUT1 0 VALUE={if(V(IN1)>{VTH}&V(IN2)>{VTH}&V(IN3)>{VTH},0,{VDD})}
R3 OUT1 OUT {{DELAY}*1E9}
C3 OUT 0 1.443n
.ENDS NAND3_SAN
*$
.SUBCKT NAND4_SAN IN1 IN2 IN3 IN4 OUT PARAMS:VDD=5 VSS=0 VTH=2.5 DELAY=1N
E3 OUT1 0 VALUE={if(V(IN1)>VTH&V(IN2)>VTH&V(IN3)>VTH&V(IN4)>VTH,0,VDD)}
R3 OUT1 OUT {{DELAY}*1E9}
C3 OUT 0 1.443n
.ENDS NAND4_SAN
*$
.SUBCKT NOR2_SAN IN1 IN2 OUT PARAMS:VDD=5 VSS=0 VTH=2.5 DELAY =1N
E1 OUT1 0 VALUE={if(V(IN1)<{VTH}&V(IN2)<{VTH},{VDD},0)}
R5 OUT1 OUT {{DELAY}*1E9}
C5 OUT 0 1.443n
.ENDS NOR2_SAN
*$
.SUBCKT NOR3_SAN IN1 IN2 IN3 OUT PARAMS:VDD=5 VSS=0 VTH=2.5 DELAY =1N
E1 OUT1 0 VALUE={if(V(IN1)<{VTH}&V(IN2)<{VTH}&V(IN3)<{VTH},{VDD},0)}
R5 OUT1 OUT {{DELAY}*1E9}
C5 OUT 0 1.443n
.ENDS NOR3_SAN
*$
.SUBCKT NOR4_SAN IN1 IN2 IN3 IN4 OUT PARAMS:VDD=5 VSS=0 VTH=2.5 DELAY=1n
E1 OUT1 0 VALUE= {if(V(IN1)<{VTH}&V(IN2)<{VTH}&V(IN3)<{VTH}&V(IN4)<{VTH},{VDD},0)}
R5 OUT1 OUT {{DELAY}*1E9}
C5 OUT 0 1n
.ENDS NOR4_SAN
*$
.SUBCKT OR2_SAN IN1 IN2 OUT PARAMS: VDD=5 VSS=0 VTH=2.5 DELAY=1N
E1 OUT1 0 VALUE={if(V(IN1)<{VTH}&V(IN2)<{VTH},{VSS},{VDD})}
R5 OUT1 OUT {{DELAY}*1E9}
C5 OUT 0 1.443n
.ENDS OR2_SAN
*$
.SUBCKT OR3_SAN IN1 IN2 IN3 OUT PARAMS:VDD=5 VSS=0 VTH=2.5 DELAY=1N
E1 OUT1 0 VALUE={if(V(IN1)<{VTH}&V(IN2)<{VTH}&V(IN3)<{VTH},0,{VDD})}
R1 OUT1 OUT {{DELAY}*1E9}
C1 OUT 0 1.443n
.ENDS OR3_SAN
*$
.SUBCKT OR4_SAN IN1 IN2 IN3 IN4 OUT PARAMS:VDD=5 VSS=0 VTH=2.5 DELAY=1N
E1 OUT1 0 VALUE={if(V(IN1)<{VTH}&V(IN2)<{VTH}&V(IN3)<{VTH}&V(IN4)<{VTH},0,{VDD})}
R1 OUT1 OUT {{DELAY}*1E9}
C1 OUT 0 1.443n
.ENDS OR4_SAN
*$
.SUBCKT XNOR2_SAN IN1 IN2 OUT PARAMS:VDD=5 VSS=0 VTH=2.5 DELAY=1N
E1 OUT1 0 VALUE={if((V(IN1)>{VTH}&V(IN2)>{VTH})|(V(IN1)<{VTH}&V(IN2)<{VTH}),{VDD},{VSS})}
R1 OUT1 OUT {{DELAY}*1E9}
C1 OUT 0 1.443n
.ENDS XNOR2_SAN
*$
.SUBCKT XOR2_SAN IN1 IN2 OUT PARAMS:VDD=5 VSS=0 VTH=2.5 DELAY=1n
E1 OUT1 0 VALUE={if((V(IN1)>{VTH}&V(IN2)>{VTH})|(V(IN1)<{VTH}&V(IN2)<{VTH}),{VDD},{VSS})}
R1 OUT1 OUT {{DELAY}*1E9}
C1 OUT 0 1.443n
.ENDS XOR2_SAN
*$
.subckt COMPHYS2_SAN  INP INM HYS VOUT ;PARAMS: VDD=5 VSS=0 VTH=2.5 DELAY=1N
E1 VOUT_PRE 0 value = {if(V(INP)>(V(INM)+V(HYS)/2),VDD,VSS)} 
R1 VOUT_PRE VOUT {{DELAY}*1E9}
C1 VOUT 0 1.443n
.ends COMPHYS2_SAN 
*$
.SUBCKT COUNT IN RST OUT PARAMS: VDD=5 VSS=0 VTH=2.5 DELAY=1N
XU4         RST RST_B INV_DELAY_SAN PARAMS: VDD={VDD} VSS={VSS} VTH={VTH} DELAY=1N
SW5         TEMP 0 RST 0  S_VSWITCH_1
SW3         OUT 0 RST 0  S_VSWITCH_2
SW1         5 4 RST_B 0  S_VSWITCH_3
C4          3 0 1N
R2          11 3 1
ECS1        11 0 VALUE = {IF(V(IN,0)>0.9,1,0)}
C1          12 0 1.443N
XU2         IN 13 INV_DELAY_SAN PARAMS: VDD={VDD} VSS={VSS} VTH={VTH} DELAY={DELAY}
XU1         13 12 NEG_EDGE AND2_SAN PARAMS: VDD={VDD} VSS={VSS} VTH={VTH} DELAY={DELAY}
R1          IN 12 20
C3          TEMP 0 1U
XU3         8 TEMP DIODE
EVCVS2      NODE1 0 TEMP 0  1
SW2         7 8 NEG_EDGE 0  S_VSWITCH_4
EVCVS3      7 0 OUT 0  1
C2          OUT 0 1U
XD1         5 OUT DIODE
EVCVS1      4 NODE1 3 0  1
.MODEL S_VSWITCH_1 VSWITCH (RON=1M ROFF=1G VON=500M VOFF=400M)
.MODEL S_VSWITCH_2 VSWITCH (RON=1M ROFF=1G VON=800M VOFF=200M)
.MODEL S_VSWITCH_3 VSWITCH (RON=1M ROFF=1G VON=500M VOFF=400M)
.MODEL S_VSWITCH_4 VSWITCH (RON=1M ROFF=1G VON=800M VOFF=200M)
.ENDS COUNT 
*$
.SUBCKT RISE_EDGE_DETECT CLK_IN EN OUT PARAMS: PULSE_WIDTH = 1N VDD =5 VSS = 0
.PARAM VTH = {({VDD} + {VSS})/2}
C2          3 0 1.443p
EBUF        4 0 VALUE = {IF(V(3,0)>{VTH},{VSS},{VDD})}
ENAND        OUT 0 VALUE = {IF(V(4,0)<{VTH}&V(5,0)<{VTH}&V(EN,0)>{VTH},{VDD},{VSS})}
ENOT        5 0 VALUE = {IF(V(CLK_IN,0)>{VTH},{VSS},{VDD})} 
R2          3 5 {PULSE_WIDTH*1E12}
.ENDS RISE_EDGE_DETECT
*$
.SUBCKT FALL_EDGE_DETECT CLK_IN EN OUT PARAMS: PULSE_WIDTH = 1p VDD =5 VSS = 0
.PARAM VTH = {({VDD} + {VSS})/2}
C2          3 0 1.443p
ENOT2        4 0 VALUE = {IF(V(3,0)>{VTH},{VSS},{VDD})}
EAND        OUT 0 VALUE = {IF(V(4,0)>{VTH}&V(5,0)>{VTH}&V(EN,0)>{VTH},{VDD},{VSS})}
ENOT        5 0 VALUE = {IF(V(CLK_IN,0)>{VTH},{VSS},{VDD})}
R2          3 5 {PULSE_WIDTH*1E12}
.ENDS FALL_EDGE_DETECT
*$
.SUBCKT COUNTER IN_CLK EN COUNT PARAMS: MAX_COUNT = 100
IS1         4 5 1
V1          4 0 {MAX_COUNT}
SW2         0 COUNT EN 0  S_VSWITCH_1
SW1         5 COUNT 6 0  S_VSWITCH_2
C1          COUNT 0 1N
.IC V(COUNT)=0 
XU2         5 4 DIODE
XU1         IN_CLK 6 RISE_EDGE_DET_SAN_0
+ ;PARAMS: VDD=5 VSS=0 T=1N
.MODEL S_VSWITCH_1 VSWITCH (RON=1G ROFF=1U VON=500M VOFF=200M)
.MODEL S_VSWITCH_2 VSWITCH (RON=1U ROFF=1G VON=500M VOFF=200M)
.ENDS COUNTER 
*$
*RISING EDGE DETECTOR
.SUBCKT RISE_EDGE_DET_SAN_0  IN EN OUT PARAMS:VDD=5 VSS=0 T=1N
.PARAM VTH={({VDD}+{VSS})/2}
XU1 IN IN2 OUT EN AND3_SAN PARAMS:VDD=5 VSS=2.5 DELAY=1p
XU2 IN OUT_IN INV_DELAY_SAN PARAMS:VDD=5 VSS=0 VTH=2.5 DELAY=1p
XU3 OUT_IN IN2 DIODE
R1 OUT_IN IN2 {{{T}*1E12}}
C1 IN2 0 1.43P
.ENDS RISE_EDGE_DET_SAN_0 
*$
.SUBCKT SR_LATCH R S Q PARAMS: VDD=5 VSS=0 DELAY=1p VTH=2.5
C_C1         0 N00080  1p   
R_R1         0 N00080  1MEG  
X_U1         N00080 N002491 DIODE 
X_U2         0 N00080 DIODE 
X_U3         N00080 Q BUF_DELAY_SAN PARAMS: VDD={VDD} VSS={VSS} DELAY={DELAY} VTH={VTH}
V_V1         N002491 0 5
G_ABMI1         N00080 0 VALUE { if(V(R)>{VTH},{VDD},if(V(S)>{VTH},-{VDD},0))    }
.ENDS SR_LATCH 
*$
.SUBCKT SR_LATCH_SHP R S Q PARAMS: VDD=5 VSS=0 DELAY=1p VTH=2.5
C_C1         0 N00080  1p   
R_R1         0 N00080  1MEG 
X_U1         N00080 N002491 DIODE 
X_U2         0 N00080 DIODE 
X_U3         N00080 Q BUF_DELAY_SAN PARAMS: VDD={VDD} VSS={VSS} DELAY={DELAY} VTH={VTH}
V_V1         N002491 0 5
G_ABMI1         N00080 0 VALUE { if(V(S)>{VTH},-{VDD},if(V(R)>{VTH},{VDD},0))    }
.ENDS SR_LATCH_SHP 
*$
*PROGRAMMABLE CURRENT MOSFET 
.SUBCKT MOS D G S
.PARAM VTH = 0.5
.PARAM K = 2.8
E1 1 0 VALUE={IF(V(S,G)>VTH,1,0)}
G1 S D VALUE = {V(1,0)*(IF(V(S,D)> (V(S,G)-VTH),(K*V(S,G)-VTH)**2,0.5*K*(V(S,G)-VTH)*V(S,D)))}
.ENDS MOS
*$
*WITH DELAY
.SUBCKT INV_1 IN OUT VDD VSS PARAMS: DELAY=1p
E1 OUT1 0 VALUE={IF(V(IN)>{(V(VDD)+V(VSS))/2},V(VSS),V(VDD))}
R1 OUT1 OUT2 {{DELAY}*1E12}
C1 OUT2 0 1.443p
E2 OUT 0 VALUE={IF(V(OUT2)>{(V(VDD)+V(VSS))/2},V(VDD),V(VSS))}
.ENDS INV_1
*************************************** DNL Addition ***********************************
*$
.SUBCKT INL_ADD OUT IN EN
E_ABM1    OUT 0 VALUE { IF(V(EN)<0.5,0,V(N421212)) }  
E_E1         N421212 0 TABLE { V(IN, 0) }  
+((0	0)
+(3.00E+01	1.53E-06)
+(1.80E+02	-7.63E-07)
+(3.40E+02	-4.20E-06)
+(5.00E+02	-6.90E-06)
+(6.30E+02	-8.81E-06)
+(8.10E+02	-1.22E-05)
+(9.50E+02	-1.53E-05)
+(1.08E+03	-1.76E-05)
+(1.23E+03	-1.95E-05)
+(1.42E+03	-2.56E-05)
+(1.58E+03	-2.53E-05)
+(3.32E+03	-1.71E-05)
+(3.48E+03	-1.66E-05)
+(3.65E+03	-2.03E-05)
+(3.79E+03	-2.22E-05)
+(3.95E+03	-1.40E-05)
+(4.13E+03	-1.11E-05)
+(4.27E+03	-7.86E-06)
+(4.48E+03	-8.62E-06)
+(4.60E+03	-9.00E-06)
+(4.71E+03	-1.03E-05)
+(4.89E+03	-1.11E-05)
+(5.09E+03	-1.15E-05)
+(5.19E+03	-1.17E-05)
+(5.32E+03	-1.24E-05)
+(5.40E+03	-1.42E-05)
+(5.57E+03	-1.48E-05)
+(5.72E+03	-1.50E-05)
+(5.83E+03	-1.51E-05)
+(5.94E+03	-1.53E-05)
+(6.11E+03	-1.46E-05)
+(6.25E+03	-1.40E-05)
+(6.42E+03	-1.40E-05)
+(6.56E+03	-1.40E-05)
+(6.69E+03	-1.42E-05)
+(6.82E+03	-1.44E-05)
+(6.94E+03	-1.44E-05)
+(7.08E+03	-1.46E-05)
+(7.20E+03	-1.50E-05)
+(7.34E+03	-1.50E-05)
+(7.43E+03	-1.51E-05)
+(7.56E+03	-1.53E-05)
+(7.67E+03	-1.53E-05)
+(7.79E+03	-1.57E-05)
+(7.91E+03	-1.57E-05)
+(8.04E+03	-1.50E-05)
+(8.18E+03	-1.42E-05)
+(8.30E+03	-1.28E-05)
+(8.43E+03	-1.26E-05)
+(8.57E+03	-1.30E-05)
+(8.69E+03	-1.32E-05)
+(8.78E+03	-1.34E-05)
+(8.85E+03	-1.38E-05)
+(8.98E+03	-1.38E-05)
+(9.03E+03	-1.38E-05)
+(9.07E+03	-1.38E-05)
+(9.12E+03	-1.38E-05)
+(9.22E+03	-1.38E-05)
+(9.27E+03	-1.36E-05)
+(9.44E+03	-1.36E-05)
+(9.53E+03	-1.36E-05)
+(9.58E+03	-1.34E-05)
+(9.65E+03	-1.34E-05)
+(9.75E+03	-1.32E-05)
+(9.82E+03	-1.32E-05)
+(9.86E+03	-1.32E-05)
+(9.92E+03	-1.32E-05)
+(1.00E+04	-1.30E-05)
+(1.01E+04	-1.20E-05)
+(1.03E+04	-1.14E-05)
+(1.04E+04	-1.22E-05)
+(1.05E+04	-1.16E-05)
+(1.06E+04	-1.18E-05)
+(1.07E+04	-1.20E-05)
+(1.08E+04	-1.18E-05)
+(1.09E+04	-1.18E-05)
+(1.10E+04	-1.18E-05)
+(1.11E+04	-1.20E-05)
+(1.12E+04	-1.18E-05)
+(1.13E+04	-1.24E-05)
+(1.14E+04	-1.24E-05)
+(1.15E+04	-1.22E-05)
+(1.16E+04	-1.16E-05)
+(1.17E+04	-1.16E-05)
+(1.18E+04	-1.16E-05)
+(1.19E+04	-1.14E-05)
+(1.20E+04	-9.16E-06)
+(1.21E+04	-8.20E-06)
+(1.22E+04	-1.91E-06)
+(1.24E+04	-1.14E-06)
+(1.25E+04	-1.14E-06)
+(1.26E+04	-1.34E-06)
+(1.28E+04	-1.72E-06)
+(1.29E+04	-2.67E-06)
+(1.30E+04	-2.48E-06)
+(1.31E+04	-2.10E-06)
+(1.32E+04	-2.10E-06)
+(1.34E+04	-2.10E-06)
+(1.35E+04	-2.10E-06)
+(1.36E+04	-2.29E-06)
+(1.37E+04	-2.10E-06)
+(1.38E+04	-2.10E-06)
+(1.39E+04	-2.10E-06)
+(1.40E+04	-1.53E-06)
+(1.41E+04	-1.72E-06)
+(1.42E+04	-1.72E-06)
+(1.43E+04	-1.53E-06)
+(1.44E+04	-1.53E-06)
+(1.45E+04	-1.72E-06)
+(1.46E+04	-2.10E-06)
+(1.47E+04	-2.29E-06)
+(1.48E+04	-2.48E-06)
+(1.49E+04	-2.48E-06)
+(1.50E+04	-3.05E-06)
+(1.51E+04	-3.05E-06)
+(1.52E+04	-3.43E-06)
+(1.53E+04	-3.43E-06)
+(1.54E+04	-3.43E-06)
+(1.56E+04	-3.43E-06)
+(1.57E+04	-3.62E-06)
+(1.58E+04	-4.20E-06)
+(1.60E+04	-4.20E-06)
+(1.62E+04	-4.39E-06)
+(1.63E+04	-3.62E-06)
+(1.64E+04	-3.24E-06)
+(1.65E+04	-3.24E-06)
+(1.67E+04	-1.72E-06)
+(1.69E+04	-1.91E-06)
+(1.71E+04	-1.91E-06)
+(1.72E+04	-9.54E-07)
+(1.74E+04	-5.72E-07)
+(1.75E+04	-5.72E-07)
+(1.76E+04	-5.72E-07)
+(1.78E+04	-5.72E-07)
+(1.79E+04	-1.91E-07)
+(1.80E+04	-9.54E-07)
+(1.81E+04	-3.43E-06)
+(1.82E+04	-4.01E-06)
+(1.83E+04	-4.01E-06)
+(1.84E+04	-4.01E-06)
+(1.85E+04	-3.62E-06)
+(1.86E+04	-3.43E-06)
+(1.87E+04	-3.62E-06)
+(1.89E+04	-3.05E-06)
+(1.91E+04	-3.24E-06)
+(1.92E+04	-3.24E-06)
+(1.93E+04	-3.62E-06)
+(1.94E+04	-3.81E-06)
+(1.95E+04	-3.24E-06)
+(1.96E+04	-3.05E-06)
+(1.97E+04	-3.24E-06)
+(1.98E+04	-3.62E-06)
+(2.00E+04	-1.14E-06)
+(2.01E+04	-5.72E-07)
+(2.02E+04	-3.81E-07)
+(2.03E+04	3.81E-07)
+(2.04E+04	3.81E-07)
+(2.05E+04	7.63E-07)
+(2.06E+04	1.72E-06)
+(2.08E+04	2.67E-06)
+(2.09E+04	3.05E-06)
+(2.11E+04	2.86E-06)
+(2.12E+04	2.67E-06)
+(2.13E+04	2.48E-06)
+(2.14E+04	2.48E-06)
+(2.15E+04	2.29E-06)
+(2.17E+04	2.29E-06)
+(2.18E+04	2.10E-06)
+(2.19E+04	2.10E-06)
+(2.20E+04	2.29E-06)
+(2.21E+04	2.29E-06)
+(2.22E+04	2.10E-06)
+(2.23E+04	2.10E-06)
+(2.24E+04	1.72E-06)
+(2.25E+04	1.72E-06)
+(2.26E+04	1.91E-06)
+(2.27E+04	2.10E-06)
+(2.28E+04	2.10E-06)
+(2.29E+04	2.29E-06)
+(2.30E+04	2.48E-06)
+(2.31E+04	2.86E-06)
+(2.32E+04	2.67E-06)
+(2.33E+04	2.48E-06)
+(2.34E+04	2.48E-06)
+(2.35E+04	2.29E-06)
+(2.36E+04	2.48E-06)
+(2.37E+04	2.48E-06)
+(2.39E+04	3.05E-06)
+(2.40E+04	2.86E-06)
+(2.42E+04	2.29E-06)
+(2.43E+04	2.48E-06)
+(2.44E+04	2.48E-06)
+(2.45E+04	2.48E-06)
+(2.46E+04	3.05E-06)
+(2.47E+04	3.24E-06)
+(2.49E+04	4.96E-06)
+(2.51E+04	5.91E-06)
+(2.52E+04	6.29E-06)
+(2.53E+04	6.29E-06)
+(2.54E+04	6.48E-06)
+(2.55E+04	7.63E-06)
+(2.56E+04	8.01E-06)
+(2.57E+04	7.06E-06)
+(2.58E+04	5.15E-06)
+(2.59E+04	4.01E-06)
+(2.60E+04	3.81E-06)
+(2.61E+04	4.01E-06)
+(2.62E+04	4.20E-06)
+(2.63E+04	4.39E-06)
+(2.64E+04	4.77E-06)
+(2.65E+04	5.72E-06)
+(2.66E+04	6.29E-06)
+(2.67E+04	6.87E-06)
+(2.68E+04	6.87E-06)
+(2.69E+04	5.34E-06)
+(2.70E+04	3.62E-06)
+(2.71E+04	4.20E-06)
+(2.72E+04	4.39E-06)
+(2.74E+04	4.39E-06)
+(2.75E+04	4.58E-06)
+(2.76E+04	4.77E-06)
+(2.77E+04	4.96E-06)
+(2.78E+04	4.96E-06)
+(2.79E+04	4.96E-06)
+(2.80E+04	4.77E-06)
+(2.81E+04	3.24E-06)
+(2.82E+04	2.29E-06)
+(2.83E+04	2.86E-06)
+(2.84E+04	3.43E-06)
+(2.85E+04	3.81E-06)
+(2.86E+04	4.77E-06)
+(2.87E+04	4.20E-06)
+(2.88E+04	6.10E-06)
+(2.89E+04	6.29E-06)
+(2.91E+04	6.10E-06)
+(2.92E+04	5.91E-06)
+(2.93E+04	4.77E-06)
+(2.94E+04	4.77E-06)
+(2.95E+04	4.77E-06)
+(2.96E+04	4.77E-06)
+(2.97E+04	4.77E-06)
+(2.98E+04	4.77E-06)
+(2.99E+04	4.20E-06)
+(3.00E+04	1.91E-06)
+(3.01E+04	1.75E-06)
+(3.03E+04	1.75E-06)
+(3.04E+04	1.79E-06)
+(3.05E+04	2.75E-06)
+(3.06E+04	2.78E-06)
+(3.07E+04	2.40E-06)
+(3.08E+04	2.59E-06)
+(3.09E+04	2.82E-06)
+(3.10E+04	4.20E-06)
+(3.11E+04	3.81E-06)
+(3.12E+04	3.81E-06)
+(3.13E+04	3.66E-06)
+(3.14E+04	3.66E-06)
+(3.15E+04	4.27E-06)
+(3.16E+04	4.27E-06)
+(3.17E+04	4.27E-06)
+(3.18E+04	4.31E-06)
+(3.19E+04	4.12E-06)
+(3.20E+04	3.74E-06)
+(3.21E+04	3.20E-06)
+(3.22E+04	3.01E-06)
+(3.23E+04	3.24E-06)
+(3.24E+04	3.43E-06)
+(3.25E+04	3.43E-06)
+(3.26E+04	4.04E-06)
+(3.27E+04	4.08E-06)
+(3.28E+04	4.08E-06)
+(3.29E+04	4.08E-06)
+(3.30E+04	4.31E-06)
+(3.31E+04	5.65E-06)
+(3.32E+04	6.64E-06)
+(3.33E+04	6.64E-06)
+(3.34E+04	6.87E-06)
+(3.35E+04	6.87E-06)
+(3.37E+04	7.67E-06)
+(3.38E+04	7.29E-06)
+(3.39E+04	7.32E-06)
+(3.40E+04	7.32E-06)
+(3.41E+04	7.13E-06)
+(3.43E+04	6.98E-06)
+(3.44E+04	7.59E-06)
+(3.45E+04	7.40E-06)
+(3.47E+04	7.06E-06)
+(3.48E+04	7.86E-06)
+(3.49E+04	8.24E-06)
+(3.50E+04	8.43E-06)
+(3.51E+04	8.47E-06)
+(3.52E+04	9.42E-06)
+(3.54E+04	1.02E-05)
+(3.55E+04	1.06E-05)
+(3.56E+04	1.12E-05)
+(3.57E+04	1.16E-05)
+(3.58E+04	1.20E-05)
+(3.60E+04	1.28E-05)
+(3.61E+04	1.19E-05)
+(3.62E+04	1.11E-05)
+(3.63E+04	9.99E-06)
+(3.64E+04	9.80E-06)
+(3.65E+04	1.00E-05)
+(3.66E+04	1.06E-05)
+(3.67E+04	1.24E-05)
+(3.69E+04	1.54E-05)
+(3.70E+04	1.70E-05)
+(3.71E+04	1.85E-05)
+(3.72E+04	1.99E-05)
+(3.74E+04	2.13E-05)
+(3.75E+04	2.32E-05)
+(3.76E+04	2.38E-05)
+(3.78E+04	2.42E-05)
+(3.79E+04	2.45E-05)
+(3.80E+04	2.48E-05)
+(3.82E+04	2.49E-05)
+(3.83E+04	2.49E-05)
+(3.84E+04	2.47E-05)
+(3.85E+04	2.51E-05)
+(3.87E+04	2.53E-05)
+(3.88E+04	2.55E-05)
+(3.89E+04	2.56E-05)
+(3.90E+04	2.50E-05)
+(3.91E+04	2.50E-05)
+(3.92E+04	2.46E-05)
+(3.93E+04	2.48E-05)
+(3.94E+04	2.46E-05)
+(3.95E+04	2.47E-05)
+(3.96E+04	2.43E-05)
+(3.97E+04	2.43E-05)
+(3.98E+04	2.43E-05)
+(3.99E+04	2.44E-05)
+(4.01E+04	2.39E-05)
+(4.02E+04	2.39E-05)
+(4.03E+04	2.39E-05)
+(4.04E+04	2.35E-05)
+(4.05E+04	2.24E-05)
+(4.07E+04	2.48E-05)
+(4.08E+04	2.85E-05)
+(4.09E+04	2.94E-05)
+(4.10E+04	3.06E-05)
+(4.11E+04	3.12E-05)
+(4.12E+04	3.14E-05)
+(4.13E+04	3.21E-05)
+(4.15E+04	3.19E-05)
+(4.16E+04	3.19E-05)
+(4.17E+04	3.23E-05)
+(4.18E+04	3.21E-05)
+(4.19E+04	3.21E-05)
+(4.21E+04	3.19E-05)
+(4.22E+04	3.23E-05)
+(4.23E+04	3.23E-05)
+(4.24E+04	3.23E-05)
+(4.25E+04	3.27E-05)
+(4.26E+04	3.27E-05)
+(4.27E+04	3.29E-05)
+(4.28E+04	3.33E-05)
+(4.30E+04	3.36E-05)
+(4.31E+04	3.42E-05)
+(4.32E+04	3.42E-05)
+(4.33E+04	3.40E-05)
+(4.34E+04	3.40E-05)
+(4.35E+04	3.57E-05)
+(4.36E+04	3.56E-05)
+(4.37E+04	3.57E-05)
+(4.38E+04	3.73E-05)
+(4.40E+04	3.73E-05)
+(4.41E+04	3.73E-05)
+(4.42E+04	3.69E-05)
+(4.44E+04	3.67E-05)
+(4.45E+04	3.56E-05)
+(4.46E+04	3.54E-05)
+(4.47E+04	3.52E-05)
+(4.48E+04	3.50E-05)
+(4.49E+04	3.48E-05)
+(4.50E+04	3.54E-05)
+(4.51E+04	3.57E-05)
+(4.52E+04	3.57E-05)
+(4.54E+04	3.57E-05)
+(4.55E+04	3.61E-05)
+(4.56E+04	3.63E-05)
+(4.57E+04	3.65E-05)
+(4.58E+04	3.67E-05)
+(4.59E+04	3.69E-05)
+(4.60E+04	3.71E-05)
+(4.61E+04	3.71E-05)
+(4.62E+04	3.71E-05)
+(4.64E+04	3.67E-05)
+(4.65E+04	3.67E-05)
+(4.66E+04	3.67E-05)
+(4.67E+04	3.73E-05)
+(4.68E+04	3.73E-05)
+(4.69E+04	3.75E-05)
+(4.71E+04	3.77E-05)
+(4.72E+04	3.84E-05)
+(4.73E+04	3.92E-05)
+(4.74E+04	3.96E-05)
+(4.75E+04	3.94E-05)
+(4.76E+04	3.94E-05)
+(4.77E+04	3.94E-05)
+(4.79E+04	3.94E-05)
+(4.80E+04	4.07E-05)
+(4.81E+04	4.38E-05)
+(4.83E+04	4.43E-05)
+(4.85E+04	4.59E-05)
+(4.86E+04	4.59E-05)
+(4.88E+04	4.57E-05)
+(4.89E+04	4.60E-05)
+(4.90E+04	4.66E-05)
+(4.91E+04	4.70E-05)
+(4.93E+04	4.70E-05)
+(4.94E+04	4.89E-05)
+(4.95E+04	4.89E-05)
+(4.96E+04	4.89E-05)
+(4.97E+04	5.03E-05)
+(4.99E+04	5.16E-05)
+(5.00E+04	5.28E-05)
+(5.01E+04	4.37E-05)
+(5.02E+04	4.37E-05)
+(5.03E+04	4.39E-05)
+(5.04E+04	4.37E-05)
+(5.05E+04	4.33E-05)
+(5.06E+04	4.35E-05)
+(5.07E+04	4.35E-05)
+(5.08E+04	4.29E-05)
+(5.09E+04	4.31E-05)
+(5.10E+04	4.29E-05)
+(5.11E+04	4.35E-05)
+(5.12E+04	4.31E-05)
+(5.13E+04	4.31E-05)
+(5.14E+04	4.27E-05)
+(5.15E+04	4.27E-05)
+(5.16E+04	4.29E-05)
+(5.17E+04	4.27E-05)
+(5.18E+04	4.25E-05)
+(5.19E+04	4.23E-05)
+(5.20E+04	4.23E-05)
+(5.21E+04	4.23E-05)
+(5.22E+04	4.23E-05)
+(5.23E+04	4.23E-05)
+(5.24E+04	4.17E-05)
+(5.25E+04	4.17E-05)
+(5.26E+04	4.17E-05)
+(5.27E+04	4.17E-05)
+(5.28E+04	4.17E-05)
+(5.29E+04	4.21E-05)
+(5.30E+04	4.21E-05)
+(5.31E+04	4.19E-05)
+(5.32E+04	4.17E-05)
+(5.33E+04	4.19E-05)
+(5.35E+04	4.19E-05)
+(5.36E+04	4.19E-05)
+(5.37E+04	4.19E-05)
+(5.38E+04	4.12E-05)
+(5.39E+04	4.12E-05)
+(5.40E+04	4.08E-05)
+(5.41E+04	4.06E-05)
+(5.42E+04	4.06E-05)
+(5.43E+04	4.04E-05)
+(5.44E+04	4.00E-05)
+(5.45E+04	3.79E-05)
+(5.47E+04	3.64E-05)
+(5.48E+04	3.51E-05)
+(5.49E+04	3.41E-05)
+(5.51E+04	3.31E-05)
+(5.52E+04	3.27E-05)
+(5.53E+04	3.25E-05)
+(5.55E+04	3.20E-05)
+(5.57E+04	3.06E-05)
+(5.58E+04	3.01E-05)
+(5.60E+04	2.95E-05)
+(5.61E+04	2.89E-05)
+(5.63E+04	2.87E-05)
+(5.64E+04	2.82E-05)
+(5.66E+04	2.80E-05)
+(5.67E+04	2.78E-05)
+(5.68E+04	2.76E-05)
+(5.70E+04	2.78E-05)
+(5.71E+04	2.76E-05)
+(5.72E+04	2.74E-05)
+(5.73E+04	2.74E-05)
+(5.74E+04	2.82E-05)
+(5.75E+04	2.85E-05)
+(5.76E+04	2.97E-05)
+(5.77E+04	2.99E-05)
+(5.78E+04	2.99E-05)
+(5.79E+04	2.95E-05)
+(5.80E+04	2.95E-05)
+(5.81E+04	3.01E-05)
+(5.82E+04	2.99E-05)
+(5.83E+04	2.95E-05)
+(5.84E+04	2.95E-05)
+(5.85E+04	2.93E-05)
+(5.86E+04	2.93E-05)
+(5.87E+04	2.93E-05)
+(5.88E+04	2.93E-05)
+(5.89E+04	2.89E-05)
+(5.90E+04	2.85E-05)
+(5.91E+04	2.78E-05)
+(5.93E+04	2.82E-05)
+(5.94E+04	2.82E-05)
+(5.95E+04	2.76E-05)
+(5.96E+04	2.55E-05)
+(5.97E+04	2.51E-05)
+(5.98E+04	2.47E-05)
+(5.99E+04	2.47E-05)
+(6.00E+04	2.32E-05)
+(6.01E+04	3.13E-05)
+(6.02E+04	3.13E-05)
+(6.03E+04	3.13E-05)
+(6.04E+04	3.13E-05)
+(6.05E+04	3.13E-05)
+(6.06E+04	3.13E-05)
+(6.07E+04	3.15E-05)
+(6.08E+04	3.15E-05)
+(6.09E+04	3.17E-05)
+(6.10E+04	3.15E-05)
+(6.11E+04	3.13E-05)
+(6.12E+04	3.09E-05)
+(6.13E+04	3.09E-05)
+(6.14E+04	3.09E-05)
+(6.15E+04	3.09E-05)
+(6.16E+04	3.05E-05)
+(6.17E+04	3.07E-05)
+(6.18E+04	3.07E-05)
+(6.19E+04	3.05E-05)
+(6.20E+04	3.03E-05)
+(6.21E+04	3.03E-05)
+(6.22E+04	3.01E-05)
+(6.23E+04	2.86E-05)
+(6.24E+04	2.72E-05)
+(6.25E+04	2.57E-05)
+(6.26E+04	2.40E-05)
+(6.28E+04	2.29E-05)
+(6.29E+04	2.20E-05)
+(6.30E+04	2.13E-05)
+(6.32E+04	2.13E-05)
+(6.33E+04	2.11E-05)
+(6.34E+04	2.09E-05)
+(6.35E+04	2.09E-05)
+(6.36E+04	2.05E-05)
+(6.37E+04	2.03E-05)
+(6.38E+04	2.03E-05)
+(6.40E+04	1.92E-05)
+(6.41E+04	1.90E-05)
+(6.43E+04	1.80E-05)
+(6.44E+04	1.80E-05)
+(6.45E+04	1.71E-05)
+(6.46E+04	1.51E-05)
+(6.47E+04	1.48E-05)
+(6.48E+04	1.42E-05)
+(6.49E+04	1.42E-05)
+(6.50E+04	1.42E-05)
+(6.51E+04	1.40E-05)
+(6.52E+04	1.38E-05)
+(6.53E+04	1.36E-05)
+(6.54E+04	1.32E-05)
+(6.55E+04	1.30E-05))
.ENDS INL_ADD
*$**********************      End        *********************$*

